
-- IMPLEMENTA��O DE UM CIRCUITO L�GICO COMBINACIONAL A PARTIR DA TABELA DA VERDADE 1 DO ARQUIVO ANEXO (COMPLEMENTO.DOC)
-- DECLARA��O DE VARI�VEL DO TIPO VETOR NA ENTIDADE PRINCIPAL

ENTITY PROJETO04 IS
PORT ( A : IN BIT_VECTOR ( 2 DOWNTO 0 ) ;
       S : OUT BIT                    ) ;
END PROJETO04 ;

ARCHITECTURE PROJ04 OF PROJETO04 IS
BEGIN

WITH A SELECT
S <= '1' WHEN "000" ,
     '0' WHEN "001" ,
     '1' WHEN "010" ,
     '1' WHEN "011" ,
     '1' WHEN "100" ,
     '0' WHEN "101" ,
     '1' WHEN "110" ,
     '0' WHEN "111" ;
     
END PROJ04 ;