
-- IMPLEMENTA��O DE UM CIRCUITO L�GICO COMBINACIONAL A PARTIR DA TABELA DA VERDADE 1 DO ARQUIVO ANEXO (COMPLEMENTO.DOC)
-- DECLARA��O DE VARI�VEL DO TIPO VETOR NA ARQUITETURA

ENTITY PROJETO03 IS
PORT ( A, B, C : IN  BIT   ;
       S       : OUT BIT ) ;
END PROJETO03 ;

ARCHITECTURE PROJ03 OF PROJETO03 IS
SIGNAL VAR01 : BIT_VECTOR ( 2 DOWNTO 0 ) ;

BEGIN
VAR01 <= A & B & C ;

WITH VAR01 SELECT
S <= '1' WHEN "000" ,
     '0' WHEN "001" ,
     '1' WHEN "010" ,
     '1' WHEN "011" ,
     '1' WHEN "100" ,
     '0' WHEN "101" ,
     '1' WHEN "110" ,
     '0' WHEN "111" ;
     
END PROJ03 ;