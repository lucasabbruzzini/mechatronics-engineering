
-- CONTADOR ASS�NCRONO CRESCENTE DE 0 A 7 (CIRCUITO 07) DO ARQUIVO ANEXO (COMPLEMENTO.DOC)

ENTITY PROJETO13 IS
PORT ( CLOCK, INICIA : IN BIT ;
	   QOUT          : BUFFER BIT_VECTOR (2 DOWNTO 0) );
END PROJETO13 ;

ARCHITECTURE PROJ13 OF PROJETO13 IS

	COMPONENT PROJETO12
	PORT (PRN, CLRN, CLKN, J, K : IN BIT;
      Q : BUFFER BIT ) ;
	END COMPONENT; 

BEGIN

FF0 : PROJETO12 PORT MAP (J => '1', K => '1', CLKN => CLOCK,   CLRN => INICIA, PRN => '1', Q => QOUT(0));
FF1 : PROJETO12 PORT MAP (J => '1', K => '1', CLKN => QOUT(0), CLRN => INICIA, PRN => '1', Q => QOUT(1));
FF2 : PROJETO12 PORT MAP (J => '1', K => '1', CLKN => QOUT(1), CLRN => INICIA, PRN => '1', Q => QOUT(2));

END PROJ13;

-- COMPONENTE: FLIP FLOP JK MESTRE ESCRAVO COM PRESET E CLEAR

ENTITY PROJETO12 IS
PORT (PRN, CLRN, CLKN, J, K : IN BIT;
      Q : BUFFER BIT ) ;
END PROJETO12 ;

ARCHITECTURE PROJ12 OF PROJETO12 IS

BEGIN

PROCESS ( PRN, CLRN, CLKN )
	BEGIN
		IF     PRN = '0' THEN Q <= '1' ;
		ELSIF CLRN = '0' THEN Q <= '0' ;
		ELSIF CLKN = '0' AND CLKN 'EVENT THEN 
			IF    J = '1' AND K = '1' THEN Q <= NOT Q ;
		    ELSIF J = '1' AND K = '0' THEN Q <= '1' ;
		    ELSIF J = '0' AND K = '1' THEN Q <= '0' ;
			END IF ;
		END IF;
	END PROCESS ;
	Q <= Q ;
END PROJ12 ;


