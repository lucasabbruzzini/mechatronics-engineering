
-- IMPLEMENTA��O DE UM MULTIPLEXADOR 4x1 CONFORME CIRCUITO 02 DO ARQUIVO ANEXO (COMPLEMENTO.DOC)
-- DECLARA��O DE VARI�VEL DO TIPO VETOR NA ENTIDADE PRINCIPAL

ENTITY PROJETO07 IS
PORT ( D0, D1, D2, D3 : IN BIT          ; 
       A : IN BIT_VECTOR ( 1 DOWNTO 0 ) ;
       S : OUT BIT                    ) ;
END PROJETO07 ;

ARCHITECTURE PROJ07 OF PROJETO07 IS
BEGIN

WITH A SELECT
S <= D0 WHEN "00" ,
     D1 WHEN "01" ,
     D2 WHEN "10" ,
     D3 WHEN "11" ;
     
END PROJ07 ;